`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:57:31 09/14/2016 
// Design Name: 
// Module Name:    transfer_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module transfer_tb;
	reg clk, reset, read, access;
	
	wire AD, CS, RD, WR;
	
	always begin
		clk <= ~clk;
		#5;
	end
	
	initial begin
		clk <= 0;
		reset <= 1;
		#40;
		reset <= 0;
		read <= 1;
		access <= 1;
		#100;
		access <= 0;
		#1000;
		read <= 0;
		access <= 1;
		#100;
		access <= 0;
		#1000;
		$stop;
	end
	
	transfer rtc(access, read, clk, reset, AD, CS, RD, WR);	
	
endmodule
